// Global nets module 

`celldefine
module cds_globals;


supply1 vdd_;

wire e4_;

wire e3_;

wire e2_;

wire e1_;

supply0 gnd_;


endmodule
`endcelldefine
